module main

struct Point {
	x int
	y int
}
